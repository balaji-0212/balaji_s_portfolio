module mul(x,y,product);
input [7:0] x,y;
output [15:0]product;

assign product=x*y;


endmodule
